`timescale 1ns/1ns
module LookupTable(addr1, addr2, addr3, addr4, mem_pipe1, mem_pipe2, mem_pipe3, mem_pipe4);
    input [3:0] addr1;
    input [3:0] addr2;
    input [3:0] addr3;
    input [3:0] addr4;
    output reg [31:0] mem_pipe1;
    output reg [31:0] mem_pipe2;
    output reg [31:0] mem_pipe3;
    output reg [31:0] mem_pipe4;

    always @(*) begin
        case (addr1)
            4'b0000: mem_pipe1= {1'b0, 31'b1111111111111111111111111111111}; // 1
            4'b0001: mem_pipe1= {2'b11, 30'b0}; // -1/2
            4'b0010: mem_pipe1= 32'b00101010101010101010101010101010;  // 0.0101010100111111111111010101010
            4'b0011: mem_pipe1= 32'b11100000000000000000000000000000;
            4'b0100: mem_pipe1= 32'b00011001100110011001100110011001;  // 0.0011001100110011001100110011011
            4'b0101: mem_pipe1= 32'b11101010101010101010101010101011;
            4'b0110: mem_pipe1= 32'b00010010010010010010010010010010; // 1/7
            4'b0111: mem_pipe1= 32'b11110000000000000000000000000000; // -1/8
            default: mem_pipe1= 32'b0;
        endcase

        case (addr2)
            4'b0000: mem_pipe2= {1'b0, 31'b1111111111111111111111111111111}; // 1
            4'b0001: mem_pipe2= {2'b11, 30'b0}; // -1/2
            4'b0010: mem_pipe2= 32'b00101010101010101010101010101010;
            4'b0011: mem_pipe2= 32'b11100000000000000000000000000000;
            4'b0100: mem_pipe2= 32'b00011001100110011001100110011001;
            4'b0101: mem_pipe2= 32'b11101010101010101010101010101011; 
            4'b0110: mem_pipe2= 32'b00010010010010010010010010010010; // 1/7
            4'b0111: mem_pipe2=  32'b11110000000000000000000000000000;// -1/8
            default: mem_pipe2= 32'b0;
        endcase

        case (addr3)
            4'b0000: mem_pipe3= {1'b0, 31'b1111111111111111111111111111111}; // 1
            4'b0001: mem_pipe3= {2'b01, 30'b0}; // -1/2
            4'b0010: mem_pipe3= 32'b00101010101010101010101010101010;
            4'b0011: mem_pipe3= 32'b11100000000000000000000000000000;
            4'b0100: mem_pipe3= 32'b00011001100110011001100110011001;
            4'b0101: mem_pipe3= 32'b11101010101010101010101010101011;
            4'b0110: mem_pipe3= 32'b00010010010010010010010010010010; // 1/7
            4'b0111: mem_pipe3=  32'b11110000000000000000000000000000;// -1/8
            default: mem_pipe3= 32'b0;
        endcase

        case (addr4)
            4'b0000: mem_pipe4= {1'b0, 31'b1111111111111111111111111111111}; // 1
            4'b0001: mem_pipe4= {2'b01, 30'b0}; // -1/2
            4'b0010: mem_pipe4= 32'b00101010101010101010101010101010;
            4'b0011: mem_pipe4= 32'b11100000000000000000000000000000;
            4'b0100: mem_pipe4= 32'b00011001100110011001100110011001;
            4'b0101: mem_pipe4= 32'b11101010101010101010101010101011;
            4'b0110: mem_pipe4= 32'b00010010010010010010010010010010; // 1/7
            4'b0111: mem_pipe4=  32'b11110000000000000000000000000000;// -1/8
            default: mem_pipe4= 32'b0;
        endcase
    end
endmodule